// 51. Explain Inline constraints using packet type and payload length example.